library verilog;
use verilog.vl_types.all;
entity tes_ps2 is
end tes_ps2;
