library verilog;
use verilog.vl_types.all;
entity test_ps2 is
end test_ps2;
